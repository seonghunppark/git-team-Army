`timescale 1ns / 1ps



module motion_display (
    input  logic                         motion_flag,
    input  logic [                  9:0] com_x,
    input  logic [                  9:0] com_y,
    input  logic                         DE,
    input  logic [                  9:0] x_pixel,
    input  logic [                  9:0] y_pixel,
    output logic [$clog2(160*120)-1 : 0] addr,
    input  logic [                 15:0] imgData,
    output logic [                  3:0] r_port,
    output logic [                  3:0] g_port,
    output logic [                  3:0] b_port
);
    logic img_display_en;
    logic [15:0] imgData_detect;

    // assign img_display_en = DE && (x_pixel < 160) && (y_pixel < 120);
    assign img_display_en = DE && (x_pixel < 320) && (y_pixel < 240);
    // assign img_display_en = DE && (x_pixel < 640) && (y_pixel < 480);
    // assign addr = img_display_en ? (160 * y_pixel + x_pixel) : 1'bz;
    // assign addr = img_display_en ? (160 * y_pixel[9:1] + x_pixel[9:1]) : 1'bz;
    assign addr = img_display_en ? (160 * y_pixel[9:1] + x_pixel[9:1]) : 1'bz;


    always_comb begin
        r_port = 0;
        g_port = 0;
        b_port = 0;
        if (img_display_en) begin
            if ((com_x - 5 < x_pixel)&&(x_pixel < com_x+5) && (com_y - 5<y_pixel)&&(y_pixel<com_y + 5)) begin
                r_port = 4'b0;
                g_port = 4'b1111;
                b_port = 4'b0;
            end else if (motion_flag) begin
                r_port = imgData[15:12] + 4'd3;
                g_port = imgData[10:7];
                b_port = imgData[4:1];
            end else begin
                r_port = imgData[15:12];
                g_port = imgData[10:7];
                b_port = imgData[4:1];
            end
        end else begin
            r_port = 0;
            g_port = 0;
            b_port = 0;
        end
    end

endmodule

module motion_coordinate (
    // global signals
    input logic clk,
    input logic reset,
    // VGA
    input logic DE,
    input logic [9:0] x_pixel,
    input logic [9:0] y_pixel,
    // internal
    input logic motion_flag,
    // output
    output logic [9:0] com_x,  // center of mass :  (x_pixel, y_pixel)
    output logic [9:0] com_y  // center of mass :  (x_pixel, y_pixel)

);

    // 핵심로직
    // compare module에서 motion flag가 들어오면
    // motion flag 뜰 때의 x_pixel과 y_pixel값을 
    // sum값에 계속 더하고
    // 이때 나누기를 하기 위해서 sum을 몇 번 더했는지 counter값을 같이 세고
    // 픽셀을 전부 세고나면 motion flag가 뜬 pixel의 중심 좌표를 계산하고
    // 그 중심 좌표값을 motion display에 보내서
    // motion display에서 해당 중심 좌표에 원을 띄우게한다.

    logic [31 : 0] sum_x_reg;
    logic [  31:0] sum_x_next;

    logic [  31:0] sum_y_reg;
    logic [  31:0] sum_y_next;

    logic [  31:0] sum_counter_next;
    logic [  31:0] sum_counter_reg;

    logic [9 : 0] com_x_reg;
    logic [9 : 0] com_x_next;

    logic [9 : 0] com_y_reg;
    logic [9 : 0] com_y_next;


    assign com_x = com_x_reg[9:0];
    assign com_y = com_y_reg[9:0];

    always_ff @(posedge clk) begin
        if (reset) begin
            sum_x_reg       <= 0;
            sum_y_reg       <= 0;
            sum_counter_reg <= 0;
            com_x_reg       <= 0;
            com_y_reg       <= 0;
        end else begin
            sum_x_reg       <= sum_x_next;
            sum_y_reg       <= sum_y_next;
            sum_counter_reg <= sum_counter_next;
            com_x_reg       <= com_x_next;
            com_y_reg       <= com_y_next;
        end
    end

    always_comb begin
        sum_counter_next = sum_counter_reg;
        sum_x_next       = sum_x_reg;
        sum_y_next       = sum_y_reg;
        com_x_next       = com_x_reg;
        com_y_next       = com_y_reg;
        // if (DE & (x_pixel <160)&(y_pixel <120)) begin
        if (DE & (x_pixel <320)&(y_pixel <240)) begin
        // if (DE & (x_pixel <640)&(y_pixel <480)) begin
            if (motion_flag) begin
                sum_x_next       = sum_x_reg + x_pixel;
                sum_y_next       = sum_y_reg + y_pixel;
                sum_counter_next = sum_counter_reg + 1;
            end
        end 

        // if ((x_pixel == 160) & (y_pixel == 120)) begin
        if ((x_pixel == 320) & (y_pixel == 240)) begin
        // if ((x_pixel == 640) & (y_pixel == 480)) begin
            sum_x_next       = 0;
            sum_y_next       = 0;
            sum_counter_next = 0;
            if (sum_counter_reg > 0) begin
                com_x_next = sum_x_reg / sum_counter_reg;
                com_y_next = sum_y_reg / sum_counter_reg;
            end
        end

    end



endmodule
